// Code your testbench here
// or browse Examples
//The purpose of this lab is to develop reset transaction, reset sequence, reset driver
//test_da_3_seq : configuring to a particular destination port using uvm_config_db
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
