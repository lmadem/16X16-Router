typedef uvm_sequencer #(packet) packet_sequencer;
