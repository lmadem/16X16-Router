// Code your testbench here
// or browse Examples
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
