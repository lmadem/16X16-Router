// Code your testbench here
// or browse Examples
//The purpose of this lab is to implement RAL configurations - Configuring the register without RAL environment
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"