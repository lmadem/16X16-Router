// Code your testbench here
// or browse Examples
//The purpose of this lab is to develop input monitor, output monitor, output agent, in-order scoreboard, and multistream scoreboard.
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
