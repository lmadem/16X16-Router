// Code your testbench here
// or browse Examples
//The purpose of this lab is to establish communication between sequence, sequencer, and driver
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
