// Code your testbench here
// or browse Examples
//The purpose of this lab is to develop sequence library, coverage component. This is a complete environment with transactions(packet, reset_packet), sequences(packet, reset), driver, reset_driver, sequencers, input agent, reset agent, output agent, coverage, scoreboard and tests
//test_seq_lib_cfg  : To configure the sequence library to execute n number of sequences
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
