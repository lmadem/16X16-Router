// Code your testbench here
// or browse Examples
//Verification of 16X16 Router - UVM 
//The purpose of this lab is to build the skeleton environment and override the base::packet class with derived::packet_da_3 class
//test_da_3_inst.sv : Overriding the base class by instance
//test_da_3_type.sv : Overriding the base class by type
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
