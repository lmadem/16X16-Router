// Code your testbench here
// or browse Examples
//The purpose of this lab is to write the driving methods(reset, main stimulus)
`include "top.sv"
`include "interface.sv"
`include "host_interface.sv"
`include "program_router_tb.sv"
